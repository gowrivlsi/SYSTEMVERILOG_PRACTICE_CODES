interface inter(input clk,rst);

 logic rd,wr;
 logic[7:0]din;
 logic full,empty;
 logic [7:0]dout;

endinterface
