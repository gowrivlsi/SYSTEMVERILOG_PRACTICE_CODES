//===================================INTERFACE DESIGN=============================
interface tlc_intf(input clk,rst);
    string Lights;
endinterface
