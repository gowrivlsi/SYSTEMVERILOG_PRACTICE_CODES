interface dff_intf(input clk,rst);
    logic [7:0]din;
    logic [7:0]q;
endinterface
