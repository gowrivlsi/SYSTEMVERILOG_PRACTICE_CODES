//=======================================DESIGN OF INTERFACE===========================
interface comp4b_intf();
    logic [3:0]a,b;
    logic g,e,l;
endinterface
