interface logic_intf(input clk,rst);
    logic a,b;
    logic and1,not1,or1,nand1,nor1,xor1,xnor1;
endinterface
