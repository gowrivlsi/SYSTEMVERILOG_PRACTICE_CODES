//=========================================DFF INTERFACE DESIIGN=================================================
interface dff8b_intf(input c,r);
    logic [7:0]d_in;
    logic [7:0]q;
endinterface
