//=========================INTERFACE ENCODER DESIGN================== 
interface enco4b_intf();
    logic [0:3]e_i;
    logic [0:1]e_y;
endinterface
