interface  half_intf();
    logic a,b;
    logic sum,carry;

    modport tb(input sum,carry,output a,b);



endinterface
