interface enco_intf;
    logic [3:0]i;
    logic [1:0]y;

    //deco output
        logic [3:0]d_o;

        
endinterface
