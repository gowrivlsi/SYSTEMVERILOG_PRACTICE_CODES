//=========================================INTERFACE CODE================================================
interface intf;
    logic [31:0]a,b;
    logic [2:0]sel;
    logic [61:0]y,A,B,C,D,G,R,T;
endinterface
